../general/fifo_v3.sv