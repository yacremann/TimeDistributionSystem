../../general/protocol/data_frames.sv