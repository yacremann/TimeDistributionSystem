../MRAM/MRAM.sv