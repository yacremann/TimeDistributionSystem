../general/watchdog/Watchdog.sv