../../general/PayloadTransmitter/PayloadTransmitter.sv