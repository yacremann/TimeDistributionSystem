../general/SlowLink/Receiver/CDR_10b_8b.sv