../../protocol/data_frames.sv