../MRAM/SPI_RW.sv