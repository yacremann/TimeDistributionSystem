../general/FrameReceiver/FrameReceiver.sv