../general/SlowLink/Receiver/AlexanderDetectorSync.sv