../general/Trigger/Trigger.sv