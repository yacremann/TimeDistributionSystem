../general/CRC/crc_calc.sv