../../PayloadTransmitter/PayloadTransmitter.sv