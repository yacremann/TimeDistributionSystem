../general/Trigger/Delay.sv