../general/Trigger/LongDivision.sv