../../CRC/crc_calc.sv