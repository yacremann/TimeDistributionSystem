../../general/FrameReceiver/FrameReceiver.sv