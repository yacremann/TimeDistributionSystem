../general/pulse_extender/pulse_extender.sv